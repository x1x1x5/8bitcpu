module overture (clk, rst, Input_1, Input_2, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Input_1;
  input  wire [0:0] Input_2;
  output  wire [7:0] Output;

  TC_Splitter8 # (.UUID(64'd3195885122167344639 ^ UUID)) Splitter8_0 (.in({{7{1'b0}}, wire_50 }), .out0(wire_8), .out1(wire_48), .out2(wire_22), .out3(wire_17), .out4(wire_25), .out5(wire_14), .out6(wire_21), .out7(wire_55));
  TC_Decoder3 # (.UUID(64'd2699913883925215058 ^ UUID)) Decoder3_1 (.dis(1'd0), .sel0(wire_8), .sel1(wire_48), .sel2(wire_22), .out0(wire_1), .out1(wire_37), .out2(wire_34), .out3(wire_15), .out4(wire_39), .out5(wire_9), .out6(wire_13), .out7());
  TC_Decoder3 # (.UUID(64'd3311212926544707724 ^ UUID)) Decoder3_2 (.dis(1'd0), .sel0(wire_17), .sel1(wire_25), .sel2(wire_14), .out0(wire_2), .out1(wire_53), .out2(wire_0), .out3(wire_16), .out4(wire_47), .out5(wire_12), .out6(wire_40), .out7());
  TC_Decoder3 # (.UUID(64'd3974024759864549773 ^ UUID)) Decoder3_3 (.dis(1'd0), .sel0(wire_21), .sel1(wire_55), .sel2(1'd0), .out0(wire_46), .out1(wire_24), .out2(wire_3), .out3(wire_27), .out4(), .out5(), .out6(), .out7());
  TC_Counter # (.UUID(64'd2242854000475277106 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_4 (.clk(clk), .rst(rst), .save(wire_26), .in(wire_7), .out(wire_32));
  TC_Switch # (.UUID(64'd4411620797192831132 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_1), .in(wire_10), .out(wire_43));
  TC_Switch # (.UUID(64'd795781106918835647 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_37), .in(wire_10), .out(wire_41));
  TC_Switch # (.UUID(64'd3355108667291252475 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_34), .in(wire_10), .out(wire_52));
  TC_Switch # (.UUID(64'd3001038835672061860 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_4), .in(wire_10), .out(wire_57));
  TC_Switch # (.UUID(64'd3118080622297509253 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_39), .in(wire_10), .out(wire_28));
  TC_Switch # (.UUID(64'd2157305596113512381 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_9), .in(wire_10), .out(wire_58));
  TC_Switch # (.UUID(64'd1667438463012334423 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_12), .in(wire_23), .out(wire_10_5));
  TC_Switch # (.UUID(64'd1147509869468458275 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_16), .in(wire_59), .out(wire_10_1));
  TC_Switch # (.UUID(64'd4465812408012960758 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_0), .in(wire_51), .out(wire_10_0));
  TC_Switch # (.UUID(64'd3460162556717909889 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_53), .in(wire_44), .out(wire_10_2));
  TC_Switch # (.UUID(64'd753724956819988128 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_2), .in(wire_29), .out(wire_10_4));
  TC_Switch # (.UUID(64'd3344862738740074333 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_13), .in(wire_10), .out(wire_54));
  TC_Switch # (.UUID(64'd3176510617450376894 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_40), .in(wire_35), .out(wire_10_6));
  TC_Switch # (.UUID(64'd1926946784219524756 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_47), .in(wire_60), .out(wire_10_3));
  TC_Switch # (.UUID(64'd4138163018043365279 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_24), .in(wire_38), .out(wire_49));
  TC_Or # (.UUID(64'd1533107826338821890 ^ UUID), .BIT_WIDTH(64'd1)) Or_20 (.in0(wire_24), .in1(wire_4), .out(wire_19));
  TC_Maker8 # (.UUID(64'd207153706724710286 ^ UUID)) Maker8_21 (.in0(wire_8), .in1(wire_48), .in2(wire_22), .in3(wire_17), .in4(wire_25), .in5(wire_14), .in6(wire_21), .in7(wire_55), .out(wire_20));
  TC_Mux # (.UUID(64'd1964629266523616625 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_22 (.sel(wire_24), .in0(wire_57), .in1(wire_49), .out(wire_45));
  TC_Switch # (.UUID(64'd99064881001667093 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_46), .in({{7{1'b0}}, wire_50 }), .out(wire_56));
  TC_Mux # (.UUID(64'd86638894695546479 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_24 (.sel(wire_42), .in0(wire_43), .in1(wire_56), .out(wire_36));
  TC_And # (.UUID(64'd2235740091360820880 ^ UUID), .BIT_WIDTH(64'd1)) And_25 (.in0(wire_3), .in1(wire_13), .out(wire_18));
  TC_And # (.UUID(64'd4504202246346605969 ^ UUID), .BIT_WIDTH(64'd1)) And_26 (.in0(wire_46), .in1(wire_46), .out(wire_42));
  TC_Or # (.UUID(64'd557051665834219798 ^ UUID), .BIT_WIDTH(64'd1)) Or_27 (.in0(wire_1), .in1(wire_46), .out(wire_11));
  TC_And # (.UUID(64'd3643539617608754151 ^ UUID), .BIT_WIDTH(64'd1)) And_28 (.in0(wire_40), .in1(wire_3), .out(wire_33_0));
  TC_Switch # (.UUID(64'd1684593356854366558 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_29 (.en(wire_27), .in(wire_30), .out(wire_26));
  TC_And # (.UUID(64'd824621369517961178 ^ UUID), .BIT_WIDTH(64'd1)) And_30 (.in0(wire_3), .in1(wire_15), .out(wire_4));
  RegisterPlus # (.UUID(64'd4067414350767443986 ^ UUID)) RegisterPlus_31 (.clk(clk), .rst(rst), .Load(wire_0), .Save_value(wire_52), .Save(wire_34), .Always_output(wire_6), .Output(wire_51));
  RegisterPlus # (.UUID(64'd573485098238337524 ^ UUID)) RegisterPlus_32 (.clk(clk), .rst(rst), .Load(wire_53), .Save_value(wire_41), .Save(wire_37), .Always_output(wire_31), .Output(wire_44));
  RegisterPlus # (.UUID(64'd1911715167693262826 ^ UUID)) RegisterPlus_33 (.clk(clk), .rst(rst), .Load(wire_2), .Save_value(wire_36), .Save(wire_11), .Always_output(wire_7), .Output(wire_29));
  RegisterPlus # (.UUID(64'd786948020129666723 ^ UUID)) RegisterPlus_34 (.clk(clk), .rst(rst), .Load(wire_16), .Save_value(wire_45), .Save(wire_19), .Always_output(wire_5), .Output(wire_59));
  RegisterPlus # (.UUID(64'd510126422459011973 ^ UUID)) RegisterPlus_35 (.clk(clk), .rst(rst), .Load(wire_47), .Save_value(wire_28), .Save(wire_39), .Always_output(), .Output(wire_60));
  RegisterPlus # (.UUID(64'd1438621956967896702 ^ UUID)) RegisterPlus_36 (.clk(clk), .rst(rst), .Load(wire_12), .Save_value(wire_58), .Save(wire_9), .Always_output(), .Output(wire_23));
  ALU # (.UUID(64'd836970191027515316 ^ UUID)) ALU_37 (.clk(clk), .rst(rst), .Instruction(wire_20), .Input_1(wire_31), .Input_2(wire_6), .Output(wire_38));
  COND # (.UUID(64'd2054271735338459541 ^ UUID)) COND_38 (.clk(clk), .rst(rst), .Condition(wire_20), .Input(wire_5), .Result(wire_30));
  TC_Switch # (.UUID(64'd2204582334536460964 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_39 (.en(wire_18), .in(wire_54), .out(Output));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_10_0;
  wire [7:0] wire_10_1;
  wire [7:0] wire_10_2;
  wire [7:0] wire_10_3;
  wire [7:0] wire_10_4;
  wire [7:0] wire_10_5;
  wire [7:0] wire_10_6;
  assign wire_10 = wire_10_0|wire_10_1|wire_10_2|wire_10_3|wire_10_4|wire_10_5|wire_10_6;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_29;
  wire [0:0] wire_30;
  wire [7:0] wire_31;
  wire [7:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_33_0;
  assign wire_33 = wire_33_0|Input_2;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  assign wire_35 = Input_1;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [7:0] wire_44;
  wire [7:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [7:0] wire_49;
  wire [0:0] wire_50;
  assign wire_50 = 0;
  wire [7:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  wire [7:0] wire_54;
  wire [0:0] wire_55;
  wire [7:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_58;
  wire [7:0] wire_59;
  wire [7:0] wire_60;

endmodule
